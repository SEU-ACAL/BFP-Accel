import "DPI-C" function void softmax_read_FP16_matrix(input bit en, input int line_num, output shortint line_data[1024]);
    
    
module softmax_input_fp16_line (
    input        en,
    input  [15:0] line_num,
    output [15:0] line_data_0,
    output [15:0] line_data_1,
    output [15:0] line_data_2,
    output [15:0] line_data_3,
    output [15:0] line_data_4,
    output [15:0] line_data_5,
    output [15:0] line_data_6,
    output [15:0] line_data_7,
    output [15:0] line_data_8,
    output [15:0] line_data_9,
    output [15:0] line_data_10,
    output [15:0] line_data_11,
    output [15:0] line_data_12,
    output [15:0] line_data_13,
    output [15:0] line_data_14,
    output [15:0] line_data_15,
    output [15:0] line_data_16,
    output [15:0] line_data_17,
    output [15:0] line_data_18,
    output [15:0] line_data_19,
    output [15:0] line_data_20,
    output [15:0] line_data_21,
    output [15:0] line_data_22,
    output [15:0] line_data_23,
    output [15:0] line_data_24,
    output [15:0] line_data_25,
    output [15:0] line_data_26,
    output [15:0] line_data_27,
    output [15:0] line_data_28,
    output [15:0] line_data_29,
    output [15:0] line_data_30,
    output [15:0] line_data_31,
    output [15:0] line_data_32,
    output [15:0] line_data_33,
    output [15:0] line_data_34,
    output [15:0] line_data_35,
    output [15:0] line_data_36,
    output [15:0] line_data_37,
    output [15:0] line_data_38,
    output [15:0] line_data_39,
    output [15:0] line_data_40,
    output [15:0] line_data_41,
    output [15:0] line_data_42,
    output [15:0] line_data_43,
    output [15:0] line_data_44,
    output [15:0] line_data_45,
    output [15:0] line_data_46,
    output [15:0] line_data_47,
    output [15:0] line_data_48,
    output [15:0] line_data_49,
    output [15:0] line_data_50,
    output [15:0] line_data_51,
    output [15:0] line_data_52,
    output [15:0] line_data_53,
    output [15:0] line_data_54,
    output [15:0] line_data_55,
    output [15:0] line_data_56,
    output [15:0] line_data_57,
    output [15:0] line_data_58,
    output [15:0] line_data_59,
    output [15:0] line_data_60,
    output [15:0] line_data_61,
    output [15:0] line_data_62,
    output [15:0] line_data_63,
    output [15:0] line_data_64,
    output [15:0] line_data_65,
    output [15:0] line_data_66,
    output [15:0] line_data_67,
    output [15:0] line_data_68,
    output [15:0] line_data_69,
    output [15:0] line_data_70,
    output [15:0] line_data_71,
    output [15:0] line_data_72,
    output [15:0] line_data_73,
    output [15:0] line_data_74,
    output [15:0] line_data_75,
    output [15:0] line_data_76,
    output [15:0] line_data_77,
    output [15:0] line_data_78,
    output [15:0] line_data_79,
    output [15:0] line_data_80,
    output [15:0] line_data_81,
    output [15:0] line_data_82,
    output [15:0] line_data_83,
    output [15:0] line_data_84,
    output [15:0] line_data_85,
    output [15:0] line_data_86,
    output [15:0] line_data_87,
    output [15:0] line_data_88,
    output [15:0] line_data_89,
    output [15:0] line_data_90,
    output [15:0] line_data_91,
    output [15:0] line_data_92,
    output [15:0] line_data_93,
    output [15:0] line_data_94,
    output [15:0] line_data_95,
    output [15:0] line_data_96,
    output [15:0] line_data_97,
    output [15:0] line_data_98,
    output [15:0] line_data_99,
    output [15:0] line_data_100,
    output [15:0] line_data_101,
    output [15:0] line_data_102,
    output [15:0] line_data_103,
    output [15:0] line_data_104,
    output [15:0] line_data_105,
    output [15:0] line_data_106,
    output [15:0] line_data_107,
    output [15:0] line_data_108,
    output [15:0] line_data_109,
    output [15:0] line_data_110,
    output [15:0] line_data_111,
    output [15:0] line_data_112,
    output [15:0] line_data_113,
    output [15:0] line_data_114,
    output [15:0] line_data_115,
    output [15:0] line_data_116,
    output [15:0] line_data_117,
    output [15:0] line_data_118,
    output [15:0] line_data_119,
    output [15:0] line_data_120,
    output [15:0] line_data_121,
    output [15:0] line_data_122,
    output [15:0] line_data_123,
    output [15:0] line_data_124,
    output [15:0] line_data_125,
    output [15:0] line_data_126,
    output [15:0] line_data_127,
    output [15:0] line_data_128,
    output [15:0] line_data_129,
    output [15:0] line_data_130,
    output [15:0] line_data_131,
    output [15:0] line_data_132,
    output [15:0] line_data_133,
    output [15:0] line_data_134,
    output [15:0] line_data_135,
    output [15:0] line_data_136,
    output [15:0] line_data_137,
    output [15:0] line_data_138,
    output [15:0] line_data_139,
    output [15:0] line_data_140,
    output [15:0] line_data_141,
    output [15:0] line_data_142,
    output [15:0] line_data_143,
    output [15:0] line_data_144,
    output [15:0] line_data_145,
    output [15:0] line_data_146,
    output [15:0] line_data_147,
    output [15:0] line_data_148,
    output [15:0] line_data_149,
    output [15:0] line_data_150,
    output [15:0] line_data_151,
    output [15:0] line_data_152,
    output [15:0] line_data_153,
    output [15:0] line_data_154,
    output [15:0] line_data_155,
    output [15:0] line_data_156,
    output [15:0] line_data_157,
    output [15:0] line_data_158,
    output [15:0] line_data_159,
    output [15:0] line_data_160,
    output [15:0] line_data_161,
    output [15:0] line_data_162,
    output [15:0] line_data_163,
    output [15:0] line_data_164,
    output [15:0] line_data_165,
    output [15:0] line_data_166,
    output [15:0] line_data_167,
    output [15:0] line_data_168,
    output [15:0] line_data_169,
    output [15:0] line_data_170,
    output [15:0] line_data_171,
    output [15:0] line_data_172,
    output [15:0] line_data_173,
    output [15:0] line_data_174,
    output [15:0] line_data_175,
    output [15:0] line_data_176,
    output [15:0] line_data_177,
    output [15:0] line_data_178,
    output [15:0] line_data_179,
    output [15:0] line_data_180,
    output [15:0] line_data_181,
    output [15:0] line_data_182,
    output [15:0] line_data_183,
    output [15:0] line_data_184,
    output [15:0] line_data_185,
    output [15:0] line_data_186,
    output [15:0] line_data_187,
    output [15:0] line_data_188,
    output [15:0] line_data_189,
    output [15:0] line_data_190,
    output [15:0] line_data_191,
    output [15:0] line_data_192,
    output [15:0] line_data_193,
    output [15:0] line_data_194,
    output [15:0] line_data_195,
    output [15:0] line_data_196,
    output [15:0] line_data_197,
    output [15:0] line_data_198,
    output [15:0] line_data_199,
    output [15:0] line_data_200,
    output [15:0] line_data_201,
    output [15:0] line_data_202,
    output [15:0] line_data_203,
    output [15:0] line_data_204,
    output [15:0] line_data_205,
    output [15:0] line_data_206,
    output [15:0] line_data_207,
    output [15:0] line_data_208,
    output [15:0] line_data_209,
    output [15:0] line_data_210,
    output [15:0] line_data_211,
    output [15:0] line_data_212,
    output [15:0] line_data_213,
    output [15:0] line_data_214,
    output [15:0] line_data_215,
    output [15:0] line_data_216,
    output [15:0] line_data_217,
    output [15:0] line_data_218,
    output [15:0] line_data_219,
    output [15:0] line_data_220,
    output [15:0] line_data_221,
    output [15:0] line_data_222,
    output [15:0] line_data_223,
    output [15:0] line_data_224,
    output [15:0] line_data_225,
    output [15:0] line_data_226,
    output [15:0] line_data_227,
    output [15:0] line_data_228,
    output [15:0] line_data_229,
    output [15:0] line_data_230,
    output [15:0] line_data_231,
    output [15:0] line_data_232,
    output [15:0] line_data_233,
    output [15:0] line_data_234,
    output [15:0] line_data_235,
    output [15:0] line_data_236,
    output [15:0] line_data_237,
    output [15:0] line_data_238,
    output [15:0] line_data_239,
    output [15:0] line_data_240,
    output [15:0] line_data_241,
    output [15:0] line_data_242,
    output [15:0] line_data_243,
    output [15:0] line_data_244,
    output [15:0] line_data_245,
    output [15:0] line_data_246,
    output [15:0] line_data_247,
    output [15:0] line_data_248,
    output [15:0] line_data_249,
    output [15:0] line_data_250,
    output [15:0] line_data_251,
    output [15:0] line_data_252,
    output [15:0] line_data_253,
    output [15:0] line_data_254,
    output [15:0] line_data_255,
    output [15:0] line_data_256,
    output [15:0] line_data_257,
    output [15:0] line_data_258,
    output [15:0] line_data_259,
    output [15:0] line_data_260,
    output [15:0] line_data_261,
    output [15:0] line_data_262,
    output [15:0] line_data_263,
    output [15:0] line_data_264,
    output [15:0] line_data_265,
    output [15:0] line_data_266,
    output [15:0] line_data_267,
    output [15:0] line_data_268,
    output [15:0] line_data_269,
    output [15:0] line_data_270,
    output [15:0] line_data_271,
    output [15:0] line_data_272,
    output [15:0] line_data_273,
    output [15:0] line_data_274,
    output [15:0] line_data_275,
    output [15:0] line_data_276,
    output [15:0] line_data_277,
    output [15:0] line_data_278,
    output [15:0] line_data_279,
    output [15:0] line_data_280,
    output [15:0] line_data_281,
    output [15:0] line_data_282,
    output [15:0] line_data_283,
    output [15:0] line_data_284,
    output [15:0] line_data_285,
    output [15:0] line_data_286,
    output [15:0] line_data_287,
    output [15:0] line_data_288,
    output [15:0] line_data_289,
    output [15:0] line_data_290,
    output [15:0] line_data_291,
    output [15:0] line_data_292,
    output [15:0] line_data_293,
    output [15:0] line_data_294,
    output [15:0] line_data_295,
    output [15:0] line_data_296,
    output [15:0] line_data_297,
    output [15:0] line_data_298,
    output [15:0] line_data_299,
    output [15:0] line_data_300,
    output [15:0] line_data_301,
    output [15:0] line_data_302,
    output [15:0] line_data_303,
    output [15:0] line_data_304,
    output [15:0] line_data_305,
    output [15:0] line_data_306,
    output [15:0] line_data_307,
    output [15:0] line_data_308,
    output [15:0] line_data_309,
    output [15:0] line_data_310,
    output [15:0] line_data_311,
    output [15:0] line_data_312,
    output [15:0] line_data_313,
    output [15:0] line_data_314,
    output [15:0] line_data_315,
    output [15:0] line_data_316,
    output [15:0] line_data_317,
    output [15:0] line_data_318,
    output [15:0] line_data_319,
    output [15:0] line_data_320,
    output [15:0] line_data_321,
    output [15:0] line_data_322,
    output [15:0] line_data_323,
    output [15:0] line_data_324,
    output [15:0] line_data_325,
    output [15:0] line_data_326,
    output [15:0] line_data_327,
    output [15:0] line_data_328,
    output [15:0] line_data_329,
    output [15:0] line_data_330,
    output [15:0] line_data_331,
    output [15:0] line_data_332,
    output [15:0] line_data_333,
    output [15:0] line_data_334,
    output [15:0] line_data_335,
    output [15:0] line_data_336,
    output [15:0] line_data_337,
    output [15:0] line_data_338,
    output [15:0] line_data_339,
    output [15:0] line_data_340,
    output [15:0] line_data_341,
    output [15:0] line_data_342,
    output [15:0] line_data_343,
    output [15:0] line_data_344,
    output [15:0] line_data_345,
    output [15:0] line_data_346,
    output [15:0] line_data_347,
    output [15:0] line_data_348,
    output [15:0] line_data_349,
    output [15:0] line_data_350,
    output [15:0] line_data_351,
    output [15:0] line_data_352,
    output [15:0] line_data_353,
    output [15:0] line_data_354,
    output [15:0] line_data_355,
    output [15:0] line_data_356,
    output [15:0] line_data_357,
    output [15:0] line_data_358,
    output [15:0] line_data_359,
    output [15:0] line_data_360,
    output [15:0] line_data_361,
    output [15:0] line_data_362,
    output [15:0] line_data_363,
    output [15:0] line_data_364,
    output [15:0] line_data_365,
    output [15:0] line_data_366,
    output [15:0] line_data_367,
    output [15:0] line_data_368,
    output [15:0] line_data_369,
    output [15:0] line_data_370,
    output [15:0] line_data_371,
    output [15:0] line_data_372,
    output [15:0] line_data_373,
    output [15:0] line_data_374,
    output [15:0] line_data_375,
    output [15:0] line_data_376,
    output [15:0] line_data_377,
    output [15:0] line_data_378,
    output [15:0] line_data_379,
    output [15:0] line_data_380,
    output [15:0] line_data_381,
    output [15:0] line_data_382,
    output [15:0] line_data_383,
    output [15:0] line_data_384,
    output [15:0] line_data_385,
    output [15:0] line_data_386,
    output [15:0] line_data_387,
    output [15:0] line_data_388,
    output [15:0] line_data_389,
    output [15:0] line_data_390,
    output [15:0] line_data_391,
    output [15:0] line_data_392,
    output [15:0] line_data_393,
    output [15:0] line_data_394,
    output [15:0] line_data_395,
    output [15:0] line_data_396,
    output [15:0] line_data_397,
    output [15:0] line_data_398,
    output [15:0] line_data_399,
    output [15:0] line_data_400,
    output [15:0] line_data_401,
    output [15:0] line_data_402,
    output [15:0] line_data_403,
    output [15:0] line_data_404,
    output [15:0] line_data_405,
    output [15:0] line_data_406,
    output [15:0] line_data_407,
    output [15:0] line_data_408,
    output [15:0] line_data_409,
    output [15:0] line_data_410,
    output [15:0] line_data_411,
    output [15:0] line_data_412,
    output [15:0] line_data_413,
    output [15:0] line_data_414,
    output [15:0] line_data_415,
    output [15:0] line_data_416,
    output [15:0] line_data_417,
    output [15:0] line_data_418,
    output [15:0] line_data_419,
    output [15:0] line_data_420,
    output [15:0] line_data_421,
    output [15:0] line_data_422,
    output [15:0] line_data_423,
    output [15:0] line_data_424,
    output [15:0] line_data_425,
    output [15:0] line_data_426,
    output [15:0] line_data_427,
    output [15:0] line_data_428,
    output [15:0] line_data_429,
    output [15:0] line_data_430,
    output [15:0] line_data_431,
    output [15:0] line_data_432,
    output [15:0] line_data_433,
    output [15:0] line_data_434,
    output [15:0] line_data_435,
    output [15:0] line_data_436,
    output [15:0] line_data_437,
    output [15:0] line_data_438,
    output [15:0] line_data_439,
    output [15:0] line_data_440,
    output [15:0] line_data_441,
    output [15:0] line_data_442,
    output [15:0] line_data_443,
    output [15:0] line_data_444,
    output [15:0] line_data_445,
    output [15:0] line_data_446,
    output [15:0] line_data_447,
    output [15:0] line_data_448,
    output [15:0] line_data_449,
    output [15:0] line_data_450,
    output [15:0] line_data_451,
    output [15:0] line_data_452,
    output [15:0] line_data_453,
    output [15:0] line_data_454,
    output [15:0] line_data_455,
    output [15:0] line_data_456,
    output [15:0] line_data_457,
    output [15:0] line_data_458,
    output [15:0] line_data_459,
    output [15:0] line_data_460,
    output [15:0] line_data_461,
    output [15:0] line_data_462,
    output [15:0] line_data_463,
    output [15:0] line_data_464,
    output [15:0] line_data_465,
    output [15:0] line_data_466,
    output [15:0] line_data_467,
    output [15:0] line_data_468,
    output [15:0] line_data_469,
    output [15:0] line_data_470,
    output [15:0] line_data_471,
    output [15:0] line_data_472,
    output [15:0] line_data_473,
    output [15:0] line_data_474,
    output [15:0] line_data_475,
    output [15:0] line_data_476,
    output [15:0] line_data_477,
    output [15:0] line_data_478,
    output [15:0] line_data_479,
    output [15:0] line_data_480,
    output [15:0] line_data_481,
    output [15:0] line_data_482,
    output [15:0] line_data_483,
    output [15:0] line_data_484,
    output [15:0] line_data_485,
    output [15:0] line_data_486,
    output [15:0] line_data_487,
    output [15:0] line_data_488,
    output [15:0] line_data_489,
    output [15:0] line_data_490,
    output [15:0] line_data_491,
    output [15:0] line_data_492,
    output [15:0] line_data_493,
    output [15:0] line_data_494,
    output [15:0] line_data_495,
    output [15:0] line_data_496,
    output [15:0] line_data_497,
    output [15:0] line_data_498,
    output [15:0] line_data_499,
    output [15:0] line_data_500,
    output [15:0] line_data_501,
    output [15:0] line_data_502,
    output [15:0] line_data_503,
    output [15:0] line_data_504,
    output [15:0] line_data_505,
    output [15:0] line_data_506,
    output [15:0] line_data_507,
    output [15:0] line_data_508,
    output [15:0] line_data_509,
    output [15:0] line_data_510,
    output [15:0] line_data_511,
    output [15:0] line_data_512,
    output [15:0] line_data_513,
    output [15:0] line_data_514,
    output [15:0] line_data_515,
    output [15:0] line_data_516,
    output [15:0] line_data_517,
    output [15:0] line_data_518,
    output [15:0] line_data_519,
    output [15:0] line_data_520,
    output [15:0] line_data_521,
    output [15:0] line_data_522,
    output [15:0] line_data_523,
    output [15:0] line_data_524,
    output [15:0] line_data_525,
    output [15:0] line_data_526,
    output [15:0] line_data_527,
    output [15:0] line_data_528,
    output [15:0] line_data_529,
    output [15:0] line_data_530,
    output [15:0] line_data_531,
    output [15:0] line_data_532,
    output [15:0] line_data_533,
    output [15:0] line_data_534,
    output [15:0] line_data_535,
    output [15:0] line_data_536,
    output [15:0] line_data_537,
    output [15:0] line_data_538,
    output [15:0] line_data_539,
    output [15:0] line_data_540,
    output [15:0] line_data_541,
    output [15:0] line_data_542,
    output [15:0] line_data_543,
    output [15:0] line_data_544,
    output [15:0] line_data_545,
    output [15:0] line_data_546,
    output [15:0] line_data_547,
    output [15:0] line_data_548,
    output [15:0] line_data_549,
    output [15:0] line_data_550,
    output [15:0] line_data_551,
    output [15:0] line_data_552,
    output [15:0] line_data_553,
    output [15:0] line_data_554,
    output [15:0] line_data_555,
    output [15:0] line_data_556,
    output [15:0] line_data_557,
    output [15:0] line_data_558,
    output [15:0] line_data_559,
    output [15:0] line_data_560,
    output [15:0] line_data_561,
    output [15:0] line_data_562,
    output [15:0] line_data_563,
    output [15:0] line_data_564,
    output [15:0] line_data_565,
    output [15:0] line_data_566,
    output [15:0] line_data_567,
    output [15:0] line_data_568,
    output [15:0] line_data_569,
    output [15:0] line_data_570,
    output [15:0] line_data_571,
    output [15:0] line_data_572,
    output [15:0] line_data_573,
    output [15:0] line_data_574,
    output [15:0] line_data_575,
    output [15:0] line_data_576,
    output [15:0] line_data_577,
    output [15:0] line_data_578,
    output [15:0] line_data_579,
    output [15:0] line_data_580,
    output [15:0] line_data_581,
    output [15:0] line_data_582,
    output [15:0] line_data_583,
    output [15:0] line_data_584,
    output [15:0] line_data_585,
    output [15:0] line_data_586,
    output [15:0] line_data_587,
    output [15:0] line_data_588,
    output [15:0] line_data_589,
    output [15:0] line_data_590,
    output [15:0] line_data_591,
    output [15:0] line_data_592,
    output [15:0] line_data_593,
    output [15:0] line_data_594,
    output [15:0] line_data_595,
    output [15:0] line_data_596,
    output [15:0] line_data_597,
    output [15:0] line_data_598,
    output [15:0] line_data_599,
    output [15:0] line_data_600,
    output [15:0] line_data_601,
    output [15:0] line_data_602,
    output [15:0] line_data_603,
    output [15:0] line_data_604,
    output [15:0] line_data_605,
    output [15:0] line_data_606,
    output [15:0] line_data_607,
    output [15:0] line_data_608,
    output [15:0] line_data_609,
    output [15:0] line_data_610,
    output [15:0] line_data_611,
    output [15:0] line_data_612,
    output [15:0] line_data_613,
    output [15:0] line_data_614,
    output [15:0] line_data_615,
    output [15:0] line_data_616,
    output [15:0] line_data_617,
    output [15:0] line_data_618,
    output [15:0] line_data_619,
    output [15:0] line_data_620,
    output [15:0] line_data_621,
    output [15:0] line_data_622,
    output [15:0] line_data_623,
    output [15:0] line_data_624,
    output [15:0] line_data_625,
    output [15:0] line_data_626,
    output [15:0] line_data_627,
    output [15:0] line_data_628,
    output [15:0] line_data_629,
    output [15:0] line_data_630,
    output [15:0] line_data_631,
    output [15:0] line_data_632,
    output [15:0] line_data_633,
    output [15:0] line_data_634,
    output [15:0] line_data_635,
    output [15:0] line_data_636,
    output [15:0] line_data_637,
    output [15:0] line_data_638,
    output [15:0] line_data_639,
    output [15:0] line_data_640,
    output [15:0] line_data_641,
    output [15:0] line_data_642,
    output [15:0] line_data_643,
    output [15:0] line_data_644,
    output [15:0] line_data_645,
    output [15:0] line_data_646,
    output [15:0] line_data_647,
    output [15:0] line_data_648,
    output [15:0] line_data_649,
    output [15:0] line_data_650,
    output [15:0] line_data_651,
    output [15:0] line_data_652,
    output [15:0] line_data_653,
    output [15:0] line_data_654,
    output [15:0] line_data_655,
    output [15:0] line_data_656,
    output [15:0] line_data_657,
    output [15:0] line_data_658,
    output [15:0] line_data_659,
    output [15:0] line_data_660,
    output [15:0] line_data_661,
    output [15:0] line_data_662,
    output [15:0] line_data_663,
    output [15:0] line_data_664,
    output [15:0] line_data_665,
    output [15:0] line_data_666,
    output [15:0] line_data_667,
    output [15:0] line_data_668,
    output [15:0] line_data_669,
    output [15:0] line_data_670,
    output [15:0] line_data_671,
    output [15:0] line_data_672,
    output [15:0] line_data_673,
    output [15:0] line_data_674,
    output [15:0] line_data_675,
    output [15:0] line_data_676,
    output [15:0] line_data_677,
    output [15:0] line_data_678,
    output [15:0] line_data_679,
    output [15:0] line_data_680,
    output [15:0] line_data_681,
    output [15:0] line_data_682,
    output [15:0] line_data_683,
    output [15:0] line_data_684,
    output [15:0] line_data_685,
    output [15:0] line_data_686,
    output [15:0] line_data_687,
    output [15:0] line_data_688,
    output [15:0] line_data_689,
    output [15:0] line_data_690,
    output [15:0] line_data_691,
    output [15:0] line_data_692,
    output [15:0] line_data_693,
    output [15:0] line_data_694,
    output [15:0] line_data_695,
    output [15:0] line_data_696,
    output [15:0] line_data_697,
    output [15:0] line_data_698,
    output [15:0] line_data_699,
    output [15:0] line_data_700,
    output [15:0] line_data_701,
    output [15:0] line_data_702,
    output [15:0] line_data_703,
    output [15:0] line_data_704,
    output [15:0] line_data_705,
    output [15:0] line_data_706,
    output [15:0] line_data_707,
    output [15:0] line_data_708,
    output [15:0] line_data_709,
    output [15:0] line_data_710,
    output [15:0] line_data_711,
    output [15:0] line_data_712,
    output [15:0] line_data_713,
    output [15:0] line_data_714,
    output [15:0] line_data_715,
    output [15:0] line_data_716,
    output [15:0] line_data_717,
    output [15:0] line_data_718,
    output [15:0] line_data_719,
    output [15:0] line_data_720,
    output [15:0] line_data_721,
    output [15:0] line_data_722,
    output [15:0] line_data_723,
    output [15:0] line_data_724,
    output [15:0] line_data_725,
    output [15:0] line_data_726,
    output [15:0] line_data_727,
    output [15:0] line_data_728,
    output [15:0] line_data_729,
    output [15:0] line_data_730,
    output [15:0] line_data_731,
    output [15:0] line_data_732,
    output [15:0] line_data_733,
    output [15:0] line_data_734,
    output [15:0] line_data_735,
    output [15:0] line_data_736,
    output [15:0] line_data_737,
    output [15:0] line_data_738,
    output [15:0] line_data_739,
    output [15:0] line_data_740,
    output [15:0] line_data_741,
    output [15:0] line_data_742,
    output [15:0] line_data_743,
    output [15:0] line_data_744,
    output [15:0] line_data_745,
    output [15:0] line_data_746,
    output [15:0] line_data_747,
    output [15:0] line_data_748,
    output [15:0] line_data_749,
    output [15:0] line_data_750,
    output [15:0] line_data_751,
    output [15:0] line_data_752,
    output [15:0] line_data_753,
    output [15:0] line_data_754,
    output [15:0] line_data_755,
    output [15:0] line_data_756,
    output [15:0] line_data_757,
    output [15:0] line_data_758,
    output [15:0] line_data_759,
    output [15:0] line_data_760,
    output [15:0] line_data_761,
    output [15:0] line_data_762,
    output [15:0] line_data_763,
    output [15:0] line_data_764,
    output [15:0] line_data_765,
    output [15:0] line_data_766,
    output [15:0] line_data_767,
    output [15:0] line_data_768,
    output [15:0] line_data_769,
    output [15:0] line_data_770,
    output [15:0] line_data_771,
    output [15:0] line_data_772,
    output [15:0] line_data_773,
    output [15:0] line_data_774,
    output [15:0] line_data_775,
    output [15:0] line_data_776,
    output [15:0] line_data_777,
    output [15:0] line_data_778,
    output [15:0] line_data_779,
    output [15:0] line_data_780,
    output [15:0] line_data_781,
    output [15:0] line_data_782,
    output [15:0] line_data_783,
    output [15:0] line_data_784,
    output [15:0] line_data_785,
    output [15:0] line_data_786,
    output [15:0] line_data_787,
    output [15:0] line_data_788,
    output [15:0] line_data_789,
    output [15:0] line_data_790,
    output [15:0] line_data_791,
    output [15:0] line_data_792,
    output [15:0] line_data_793,
    output [15:0] line_data_794,
    output [15:0] line_data_795,
    output [15:0] line_data_796,
    output [15:0] line_data_797,
    output [15:0] line_data_798,
    output [15:0] line_data_799,
    output [15:0] line_data_800,
    output [15:0] line_data_801,
    output [15:0] line_data_802,
    output [15:0] line_data_803,
    output [15:0] line_data_804,
    output [15:0] line_data_805,
    output [15:0] line_data_806,
    output [15:0] line_data_807,
    output [15:0] line_data_808,
    output [15:0] line_data_809,
    output [15:0] line_data_810,
    output [15:0] line_data_811,
    output [15:0] line_data_812,
    output [15:0] line_data_813,
    output [15:0] line_data_814,
    output [15:0] line_data_815,
    output [15:0] line_data_816,
    output [15:0] line_data_817,
    output [15:0] line_data_818,
    output [15:0] line_data_819,
    output [15:0] line_data_820,
    output [15:0] line_data_821,
    output [15:0] line_data_822,
    output [15:0] line_data_823,
    output [15:0] line_data_824,
    output [15:0] line_data_825,
    output [15:0] line_data_826,
    output [15:0] line_data_827,
    output [15:0] line_data_828,
    output [15:0] line_data_829,
    output [15:0] line_data_830,
    output [15:0] line_data_831,
    output [15:0] line_data_832,
    output [15:0] line_data_833,
    output [15:0] line_data_834,
    output [15:0] line_data_835,
    output [15:0] line_data_836,
    output [15:0] line_data_837,
    output [15:0] line_data_838,
    output [15:0] line_data_839,
    output [15:0] line_data_840,
    output [15:0] line_data_841,
    output [15:0] line_data_842,
    output [15:0] line_data_843,
    output [15:0] line_data_844,
    output [15:0] line_data_845,
    output [15:0] line_data_846,
    output [15:0] line_data_847,
    output [15:0] line_data_848,
    output [15:0] line_data_849,
    output [15:0] line_data_850,
    output [15:0] line_data_851,
    output [15:0] line_data_852,
    output [15:0] line_data_853,
    output [15:0] line_data_854,
    output [15:0] line_data_855,
    output [15:0] line_data_856,
    output [15:0] line_data_857,
    output [15:0] line_data_858,
    output [15:0] line_data_859,
    output [15:0] line_data_860,
    output [15:0] line_data_861,
    output [15:0] line_data_862,
    output [15:0] line_data_863,
    output [15:0] line_data_864,
    output [15:0] line_data_865,
    output [15:0] line_data_866,
    output [15:0] line_data_867,
    output [15:0] line_data_868,
    output [15:0] line_data_869,
    output [15:0] line_data_870,
    output [15:0] line_data_871,
    output [15:0] line_data_872,
    output [15:0] line_data_873,
    output [15:0] line_data_874,
    output [15:0] line_data_875,
    output [15:0] line_data_876,
    output [15:0] line_data_877,
    output [15:0] line_data_878,
    output [15:0] line_data_879,
    output [15:0] line_data_880,
    output [15:0] line_data_881,
    output [15:0] line_data_882,
    output [15:0] line_data_883,
    output [15:0] line_data_884,
    output [15:0] line_data_885,
    output [15:0] line_data_886,
    output [15:0] line_data_887,
    output [15:0] line_data_888,
    output [15:0] line_data_889,
    output [15:0] line_data_890,
    output [15:0] line_data_891,
    output [15:0] line_data_892,
    output [15:0] line_data_893,
    output [15:0] line_data_894,
    output [15:0] line_data_895,
    output [15:0] line_data_896,
    output [15:0] line_data_897,
    output [15:0] line_data_898,
    output [15:0] line_data_899,
    output [15:0] line_data_900,
    output [15:0] line_data_901,
    output [15:0] line_data_902,
    output [15:0] line_data_903,
    output [15:0] line_data_904,
    output [15:0] line_data_905,
    output [15:0] line_data_906,
    output [15:0] line_data_907,
    output [15:0] line_data_908,
    output [15:0] line_data_909,
    output [15:0] line_data_910,
    output [15:0] line_data_911,
    output [15:0] line_data_912,
    output [15:0] line_data_913,
    output [15:0] line_data_914,
    output [15:0] line_data_915,
    output [15:0] line_data_916,
    output [15:0] line_data_917,
    output [15:0] line_data_918,
    output [15:0] line_data_919,
    output [15:0] line_data_920,
    output [15:0] line_data_921,
    output [15:0] line_data_922,
    output [15:0] line_data_923,
    output [15:0] line_data_924,
    output [15:0] line_data_925,
    output [15:0] line_data_926,
    output [15:0] line_data_927,
    output [15:0] line_data_928,
    output [15:0] line_data_929,
    output [15:0] line_data_930,
    output [15:0] line_data_931,
    output [15:0] line_data_932,
    output [15:0] line_data_933,
    output [15:0] line_data_934,
    output [15:0] line_data_935,
    output [15:0] line_data_936,
    output [15:0] line_data_937,
    output [15:0] line_data_938,
    output [15:0] line_data_939,
    output [15:0] line_data_940,
    output [15:0] line_data_941,
    output [15:0] line_data_942,
    output [15:0] line_data_943,
    output [15:0] line_data_944,
    output [15:0] line_data_945,
    output [15:0] line_data_946,
    output [15:0] line_data_947,
    output [15:0] line_data_948,
    output [15:0] line_data_949,
    output [15:0] line_data_950,
    output [15:0] line_data_951,
    output [15:0] line_data_952,
    output [15:0] line_data_953,
    output [15:0] line_data_954,
    output [15:0] line_data_955,
    output [15:0] line_data_956,
    output [15:0] line_data_957,
    output [15:0] line_data_958,
    output [15:0] line_data_959,
    output [15:0] line_data_960,
    output [15:0] line_data_961,
    output [15:0] line_data_962,
    output [15:0] line_data_963,
    output [15:0] line_data_964,
    output [15:0] line_data_965,
    output [15:0] line_data_966,
    output [15:0] line_data_967,
    output [15:0] line_data_968,
    output [15:0] line_data_969,
    output [15:0] line_data_970,
    output [15:0] line_data_971,
    output [15:0] line_data_972,
    output [15:0] line_data_973,
    output [15:0] line_data_974,
    output [15:0] line_data_975,
    output [15:0] line_data_976,
    output [15:0] line_data_977,
    output [15:0] line_data_978,
    output [15:0] line_data_979,
    output [15:0] line_data_980,
    output [15:0] line_data_981,
    output [15:0] line_data_982,
    output [15:0] line_data_983,
    output [15:0] line_data_984,
    output [15:0] line_data_985,
    output [15:0] line_data_986,
    output [15:0] line_data_987,
    output [15:0] line_data_988,
    output [15:0] line_data_989,
    output [15:0] line_data_990,
    output [15:0] line_data_991,
    output [15:0] line_data_992,
    output [15:0] line_data_993,
    output [15:0] line_data_994,
    output [15:0] line_data_995,
    output [15:0] line_data_996,
    output [15:0] line_data_997,
    output [15:0] line_data_998,
    output [15:0] line_data_999,
    output [15:0] line_data_1000,
    output [15:0] line_data_1001,
    output [15:0] line_data_1002,
    output [15:0] line_data_1003,
    output [15:0] line_data_1004,
    output [15:0] line_data_1005,
    output [15:0] line_data_1006,
    output [15:0] line_data_1007,
    output [15:0] line_data_1008,
    output [15:0] line_data_1009,
    output [15:0] line_data_1010,
    output [15:0] line_data_1011,
    output [15:0] line_data_1012,
    output [15:0] line_data_1013,
    output [15:0] line_data_1014,
    output [15:0] line_data_1015,
    output [15:0] line_data_1016,
    output [15:0] line_data_1017,
    output [15:0] line_data_1018,
    output [15:0] line_data_1019,
    output [15:0] line_data_1020,
    output [15:0] line_data_1021,
    output [15:0] line_data_1022,
    output [15:0] line_data_1023
    );
       shortint line_data[1024];
    
       assign line_data_0 = line_data[0];
    assign line_data_1 = line_data[1];
    assign line_data_2 = line_data[2];
    assign line_data_3 = line_data[3];
    assign line_data_4 = line_data[4];
    assign line_data_5 = line_data[5];
    assign line_data_6 = line_data[6];
    assign line_data_7 = line_data[7];
    assign line_data_8 = line_data[8];
    assign line_data_9 = line_data[9];
    assign line_data_10 = line_data[10];
    assign line_data_11 = line_data[11];
    assign line_data_12 = line_data[12];
    assign line_data_13 = line_data[13];
    assign line_data_14 = line_data[14];
    assign line_data_15 = line_data[15];
    assign line_data_16 = line_data[16];
    assign line_data_17 = line_data[17];
    assign line_data_18 = line_data[18];
    assign line_data_19 = line_data[19];
    assign line_data_20 = line_data[20];
    assign line_data_21 = line_data[21];
    assign line_data_22 = line_data[22];
    assign line_data_23 = line_data[23];
    assign line_data_24 = line_data[24];
    assign line_data_25 = line_data[25];
    assign line_data_26 = line_data[26];
    assign line_data_27 = line_data[27];
    assign line_data_28 = line_data[28];
    assign line_data_29 = line_data[29];
    assign line_data_30 = line_data[30];
    assign line_data_31 = line_data[31];
    assign line_data_32 = line_data[32];
    assign line_data_33 = line_data[33];
    assign line_data_34 = line_data[34];
    assign line_data_35 = line_data[35];
    assign line_data_36 = line_data[36];
    assign line_data_37 = line_data[37];
    assign line_data_38 = line_data[38];
    assign line_data_39 = line_data[39];
    assign line_data_40 = line_data[40];
    assign line_data_41 = line_data[41];
    assign line_data_42 = line_data[42];
    assign line_data_43 = line_data[43];
    assign line_data_44 = line_data[44];
    assign line_data_45 = line_data[45];
    assign line_data_46 = line_data[46];
    assign line_data_47 = line_data[47];
    assign line_data_48 = line_data[48];
    assign line_data_49 = line_data[49];
    assign line_data_50 = line_data[50];
    assign line_data_51 = line_data[51];
    assign line_data_52 = line_data[52];
    assign line_data_53 = line_data[53];
    assign line_data_54 = line_data[54];
    assign line_data_55 = line_data[55];
    assign line_data_56 = line_data[56];
    assign line_data_57 = line_data[57];
    assign line_data_58 = line_data[58];
    assign line_data_59 = line_data[59];
    assign line_data_60 = line_data[60];
    assign line_data_61 = line_data[61];
    assign line_data_62 = line_data[62];
    assign line_data_63 = line_data[63];
    assign line_data_64 = line_data[64];
    assign line_data_65 = line_data[65];
    assign line_data_66 = line_data[66];
    assign line_data_67 = line_data[67];
    assign line_data_68 = line_data[68];
    assign line_data_69 = line_data[69];
    assign line_data_70 = line_data[70];
    assign line_data_71 = line_data[71];
    assign line_data_72 = line_data[72];
    assign line_data_73 = line_data[73];
    assign line_data_74 = line_data[74];
    assign line_data_75 = line_data[75];
    assign line_data_76 = line_data[76];
    assign line_data_77 = line_data[77];
    assign line_data_78 = line_data[78];
    assign line_data_79 = line_data[79];
    assign line_data_80 = line_data[80];
    assign line_data_81 = line_data[81];
    assign line_data_82 = line_data[82];
    assign line_data_83 = line_data[83];
    assign line_data_84 = line_data[84];
    assign line_data_85 = line_data[85];
    assign line_data_86 = line_data[86];
    assign line_data_87 = line_data[87];
    assign line_data_88 = line_data[88];
    assign line_data_89 = line_data[89];
    assign line_data_90 = line_data[90];
    assign line_data_91 = line_data[91];
    assign line_data_92 = line_data[92];
    assign line_data_93 = line_data[93];
    assign line_data_94 = line_data[94];
    assign line_data_95 = line_data[95];
    assign line_data_96 = line_data[96];
    assign line_data_97 = line_data[97];
    assign line_data_98 = line_data[98];
    assign line_data_99 = line_data[99];
    assign line_data_100 = line_data[100];
    assign line_data_101 = line_data[101];
    assign line_data_102 = line_data[102];
    assign line_data_103 = line_data[103];
    assign line_data_104 = line_data[104];
    assign line_data_105 = line_data[105];
    assign line_data_106 = line_data[106];
    assign line_data_107 = line_data[107];
    assign line_data_108 = line_data[108];
    assign line_data_109 = line_data[109];
    assign line_data_110 = line_data[110];
    assign line_data_111 = line_data[111];
    assign line_data_112 = line_data[112];
    assign line_data_113 = line_data[113];
    assign line_data_114 = line_data[114];
    assign line_data_115 = line_data[115];
    assign line_data_116 = line_data[116];
    assign line_data_117 = line_data[117];
    assign line_data_118 = line_data[118];
    assign line_data_119 = line_data[119];
    assign line_data_120 = line_data[120];
    assign line_data_121 = line_data[121];
    assign line_data_122 = line_data[122];
    assign line_data_123 = line_data[123];
    assign line_data_124 = line_data[124];
    assign line_data_125 = line_data[125];
    assign line_data_126 = line_data[126];
    assign line_data_127 = line_data[127];
    assign line_data_128 = line_data[128];
    assign line_data_129 = line_data[129];
    assign line_data_130 = line_data[130];
    assign line_data_131 = line_data[131];
    assign line_data_132 = line_data[132];
    assign line_data_133 = line_data[133];
    assign line_data_134 = line_data[134];
    assign line_data_135 = line_data[135];
    assign line_data_136 = line_data[136];
    assign line_data_137 = line_data[137];
    assign line_data_138 = line_data[138];
    assign line_data_139 = line_data[139];
    assign line_data_140 = line_data[140];
    assign line_data_141 = line_data[141];
    assign line_data_142 = line_data[142];
    assign line_data_143 = line_data[143];
    assign line_data_144 = line_data[144];
    assign line_data_145 = line_data[145];
    assign line_data_146 = line_data[146];
    assign line_data_147 = line_data[147];
    assign line_data_148 = line_data[148];
    assign line_data_149 = line_data[149];
    assign line_data_150 = line_data[150];
    assign line_data_151 = line_data[151];
    assign line_data_152 = line_data[152];
    assign line_data_153 = line_data[153];
    assign line_data_154 = line_data[154];
    assign line_data_155 = line_data[155];
    assign line_data_156 = line_data[156];
    assign line_data_157 = line_data[157];
    assign line_data_158 = line_data[158];
    assign line_data_159 = line_data[159];
    assign line_data_160 = line_data[160];
    assign line_data_161 = line_data[161];
    assign line_data_162 = line_data[162];
    assign line_data_163 = line_data[163];
    assign line_data_164 = line_data[164];
    assign line_data_165 = line_data[165];
    assign line_data_166 = line_data[166];
    assign line_data_167 = line_data[167];
    assign line_data_168 = line_data[168];
    assign line_data_169 = line_data[169];
    assign line_data_170 = line_data[170];
    assign line_data_171 = line_data[171];
    assign line_data_172 = line_data[172];
    assign line_data_173 = line_data[173];
    assign line_data_174 = line_data[174];
    assign line_data_175 = line_data[175];
    assign line_data_176 = line_data[176];
    assign line_data_177 = line_data[177];
    assign line_data_178 = line_data[178];
    assign line_data_179 = line_data[179];
    assign line_data_180 = line_data[180];
    assign line_data_181 = line_data[181];
    assign line_data_182 = line_data[182];
    assign line_data_183 = line_data[183];
    assign line_data_184 = line_data[184];
    assign line_data_185 = line_data[185];
    assign line_data_186 = line_data[186];
    assign line_data_187 = line_data[187];
    assign line_data_188 = line_data[188];
    assign line_data_189 = line_data[189];
    assign line_data_190 = line_data[190];
    assign line_data_191 = line_data[191];
    assign line_data_192 = line_data[192];
    assign line_data_193 = line_data[193];
    assign line_data_194 = line_data[194];
    assign line_data_195 = line_data[195];
    assign line_data_196 = line_data[196];
    assign line_data_197 = line_data[197];
    assign line_data_198 = line_data[198];
    assign line_data_199 = line_data[199];
    assign line_data_200 = line_data[200];
    assign line_data_201 = line_data[201];
    assign line_data_202 = line_data[202];
    assign line_data_203 = line_data[203];
    assign line_data_204 = line_data[204];
    assign line_data_205 = line_data[205];
    assign line_data_206 = line_data[206];
    assign line_data_207 = line_data[207];
    assign line_data_208 = line_data[208];
    assign line_data_209 = line_data[209];
    assign line_data_210 = line_data[210];
    assign line_data_211 = line_data[211];
    assign line_data_212 = line_data[212];
    assign line_data_213 = line_data[213];
    assign line_data_214 = line_data[214];
    assign line_data_215 = line_data[215];
    assign line_data_216 = line_data[216];
    assign line_data_217 = line_data[217];
    assign line_data_218 = line_data[218];
    assign line_data_219 = line_data[219];
    assign line_data_220 = line_data[220];
    assign line_data_221 = line_data[221];
    assign line_data_222 = line_data[222];
    assign line_data_223 = line_data[223];
    assign line_data_224 = line_data[224];
    assign line_data_225 = line_data[225];
    assign line_data_226 = line_data[226];
    assign line_data_227 = line_data[227];
    assign line_data_228 = line_data[228];
    assign line_data_229 = line_data[229];
    assign line_data_230 = line_data[230];
    assign line_data_231 = line_data[231];
    assign line_data_232 = line_data[232];
    assign line_data_233 = line_data[233];
    assign line_data_234 = line_data[234];
    assign line_data_235 = line_data[235];
    assign line_data_236 = line_data[236];
    assign line_data_237 = line_data[237];
    assign line_data_238 = line_data[238];
    assign line_data_239 = line_data[239];
    assign line_data_240 = line_data[240];
    assign line_data_241 = line_data[241];
    assign line_data_242 = line_data[242];
    assign line_data_243 = line_data[243];
    assign line_data_244 = line_data[244];
    assign line_data_245 = line_data[245];
    assign line_data_246 = line_data[246];
    assign line_data_247 = line_data[247];
    assign line_data_248 = line_data[248];
    assign line_data_249 = line_data[249];
    assign line_data_250 = line_data[250];
    assign line_data_251 = line_data[251];
    assign line_data_252 = line_data[252];
    assign line_data_253 = line_data[253];
    assign line_data_254 = line_data[254];
    assign line_data_255 = line_data[255];
    assign line_data_256 = line_data[256];
    assign line_data_257 = line_data[257];
    assign line_data_258 = line_data[258];
    assign line_data_259 = line_data[259];
    assign line_data_260 = line_data[260];
    assign line_data_261 = line_data[261];
    assign line_data_262 = line_data[262];
    assign line_data_263 = line_data[263];
    assign line_data_264 = line_data[264];
    assign line_data_265 = line_data[265];
    assign line_data_266 = line_data[266];
    assign line_data_267 = line_data[267];
    assign line_data_268 = line_data[268];
    assign line_data_269 = line_data[269];
    assign line_data_270 = line_data[270];
    assign line_data_271 = line_data[271];
    assign line_data_272 = line_data[272];
    assign line_data_273 = line_data[273];
    assign line_data_274 = line_data[274];
    assign line_data_275 = line_data[275];
    assign line_data_276 = line_data[276];
    assign line_data_277 = line_data[277];
    assign line_data_278 = line_data[278];
    assign line_data_279 = line_data[279];
    assign line_data_280 = line_data[280];
    assign line_data_281 = line_data[281];
    assign line_data_282 = line_data[282];
    assign line_data_283 = line_data[283];
    assign line_data_284 = line_data[284];
    assign line_data_285 = line_data[285];
    assign line_data_286 = line_data[286];
    assign line_data_287 = line_data[287];
    assign line_data_288 = line_data[288];
    assign line_data_289 = line_data[289];
    assign line_data_290 = line_data[290];
    assign line_data_291 = line_data[291];
    assign line_data_292 = line_data[292];
    assign line_data_293 = line_data[293];
    assign line_data_294 = line_data[294];
    assign line_data_295 = line_data[295];
    assign line_data_296 = line_data[296];
    assign line_data_297 = line_data[297];
    assign line_data_298 = line_data[298];
    assign line_data_299 = line_data[299];
    assign line_data_300 = line_data[300];
    assign line_data_301 = line_data[301];
    assign line_data_302 = line_data[302];
    assign line_data_303 = line_data[303];
    assign line_data_304 = line_data[304];
    assign line_data_305 = line_data[305];
    assign line_data_306 = line_data[306];
    assign line_data_307 = line_data[307];
    assign line_data_308 = line_data[308];
    assign line_data_309 = line_data[309];
    assign line_data_310 = line_data[310];
    assign line_data_311 = line_data[311];
    assign line_data_312 = line_data[312];
    assign line_data_313 = line_data[313];
    assign line_data_314 = line_data[314];
    assign line_data_315 = line_data[315];
    assign line_data_316 = line_data[316];
    assign line_data_317 = line_data[317];
    assign line_data_318 = line_data[318];
    assign line_data_319 = line_data[319];
    assign line_data_320 = line_data[320];
    assign line_data_321 = line_data[321];
    assign line_data_322 = line_data[322];
    assign line_data_323 = line_data[323];
    assign line_data_324 = line_data[324];
    assign line_data_325 = line_data[325];
    assign line_data_326 = line_data[326];
    assign line_data_327 = line_data[327];
    assign line_data_328 = line_data[328];
    assign line_data_329 = line_data[329];
    assign line_data_330 = line_data[330];
    assign line_data_331 = line_data[331];
    assign line_data_332 = line_data[332];
    assign line_data_333 = line_data[333];
    assign line_data_334 = line_data[334];
    assign line_data_335 = line_data[335];
    assign line_data_336 = line_data[336];
    assign line_data_337 = line_data[337];
    assign line_data_338 = line_data[338];
    assign line_data_339 = line_data[339];
    assign line_data_340 = line_data[340];
    assign line_data_341 = line_data[341];
    assign line_data_342 = line_data[342];
    assign line_data_343 = line_data[343];
    assign line_data_344 = line_data[344];
    assign line_data_345 = line_data[345];
    assign line_data_346 = line_data[346];
    assign line_data_347 = line_data[347];
    assign line_data_348 = line_data[348];
    assign line_data_349 = line_data[349];
    assign line_data_350 = line_data[350];
    assign line_data_351 = line_data[351];
    assign line_data_352 = line_data[352];
    assign line_data_353 = line_data[353];
    assign line_data_354 = line_data[354];
    assign line_data_355 = line_data[355];
    assign line_data_356 = line_data[356];
    assign line_data_357 = line_data[357];
    assign line_data_358 = line_data[358];
    assign line_data_359 = line_data[359];
    assign line_data_360 = line_data[360];
    assign line_data_361 = line_data[361];
    assign line_data_362 = line_data[362];
    assign line_data_363 = line_data[363];
    assign line_data_364 = line_data[364];
    assign line_data_365 = line_data[365];
    assign line_data_366 = line_data[366];
    assign line_data_367 = line_data[367];
    assign line_data_368 = line_data[368];
    assign line_data_369 = line_data[369];
    assign line_data_370 = line_data[370];
    assign line_data_371 = line_data[371];
    assign line_data_372 = line_data[372];
    assign line_data_373 = line_data[373];
    assign line_data_374 = line_data[374];
    assign line_data_375 = line_data[375];
    assign line_data_376 = line_data[376];
    assign line_data_377 = line_data[377];
    assign line_data_378 = line_data[378];
    assign line_data_379 = line_data[379];
    assign line_data_380 = line_data[380];
    assign line_data_381 = line_data[381];
    assign line_data_382 = line_data[382];
    assign line_data_383 = line_data[383];
    assign line_data_384 = line_data[384];
    assign line_data_385 = line_data[385];
    assign line_data_386 = line_data[386];
    assign line_data_387 = line_data[387];
    assign line_data_388 = line_data[388];
    assign line_data_389 = line_data[389];
    assign line_data_390 = line_data[390];
    assign line_data_391 = line_data[391];
    assign line_data_392 = line_data[392];
    assign line_data_393 = line_data[393];
    assign line_data_394 = line_data[394];
    assign line_data_395 = line_data[395];
    assign line_data_396 = line_data[396];
    assign line_data_397 = line_data[397];
    assign line_data_398 = line_data[398];
    assign line_data_399 = line_data[399];
    assign line_data_400 = line_data[400];
    assign line_data_401 = line_data[401];
    assign line_data_402 = line_data[402];
    assign line_data_403 = line_data[403];
    assign line_data_404 = line_data[404];
    assign line_data_405 = line_data[405];
    assign line_data_406 = line_data[406];
    assign line_data_407 = line_data[407];
    assign line_data_408 = line_data[408];
    assign line_data_409 = line_data[409];
    assign line_data_410 = line_data[410];
    assign line_data_411 = line_data[411];
    assign line_data_412 = line_data[412];
    assign line_data_413 = line_data[413];
    assign line_data_414 = line_data[414];
    assign line_data_415 = line_data[415];
    assign line_data_416 = line_data[416];
    assign line_data_417 = line_data[417];
    assign line_data_418 = line_data[418];
    assign line_data_419 = line_data[419];
    assign line_data_420 = line_data[420];
    assign line_data_421 = line_data[421];
    assign line_data_422 = line_data[422];
    assign line_data_423 = line_data[423];
    assign line_data_424 = line_data[424];
    assign line_data_425 = line_data[425];
    assign line_data_426 = line_data[426];
    assign line_data_427 = line_data[427];
    assign line_data_428 = line_data[428];
    assign line_data_429 = line_data[429];
    assign line_data_430 = line_data[430];
    assign line_data_431 = line_data[431];
    assign line_data_432 = line_data[432];
    assign line_data_433 = line_data[433];
    assign line_data_434 = line_data[434];
    assign line_data_435 = line_data[435];
    assign line_data_436 = line_data[436];
    assign line_data_437 = line_data[437];
    assign line_data_438 = line_data[438];
    assign line_data_439 = line_data[439];
    assign line_data_440 = line_data[440];
    assign line_data_441 = line_data[441];
    assign line_data_442 = line_data[442];
    assign line_data_443 = line_data[443];
    assign line_data_444 = line_data[444];
    assign line_data_445 = line_data[445];
    assign line_data_446 = line_data[446];
    assign line_data_447 = line_data[447];
    assign line_data_448 = line_data[448];
    assign line_data_449 = line_data[449];
    assign line_data_450 = line_data[450];
    assign line_data_451 = line_data[451];
    assign line_data_452 = line_data[452];
    assign line_data_453 = line_data[453];
    assign line_data_454 = line_data[454];
    assign line_data_455 = line_data[455];
    assign line_data_456 = line_data[456];
    assign line_data_457 = line_data[457];
    assign line_data_458 = line_data[458];
    assign line_data_459 = line_data[459];
    assign line_data_460 = line_data[460];
    assign line_data_461 = line_data[461];
    assign line_data_462 = line_data[462];
    assign line_data_463 = line_data[463];
    assign line_data_464 = line_data[464];
    assign line_data_465 = line_data[465];
    assign line_data_466 = line_data[466];
    assign line_data_467 = line_data[467];
    assign line_data_468 = line_data[468];
    assign line_data_469 = line_data[469];
    assign line_data_470 = line_data[470];
    assign line_data_471 = line_data[471];
    assign line_data_472 = line_data[472];
    assign line_data_473 = line_data[473];
    assign line_data_474 = line_data[474];
    assign line_data_475 = line_data[475];
    assign line_data_476 = line_data[476];
    assign line_data_477 = line_data[477];
    assign line_data_478 = line_data[478];
    assign line_data_479 = line_data[479];
    assign line_data_480 = line_data[480];
    assign line_data_481 = line_data[481];
    assign line_data_482 = line_data[482];
    assign line_data_483 = line_data[483];
    assign line_data_484 = line_data[484];
    assign line_data_485 = line_data[485];
    assign line_data_486 = line_data[486];
    assign line_data_487 = line_data[487];
    assign line_data_488 = line_data[488];
    assign line_data_489 = line_data[489];
    assign line_data_490 = line_data[490];
    assign line_data_491 = line_data[491];
    assign line_data_492 = line_data[492];
    assign line_data_493 = line_data[493];
    assign line_data_494 = line_data[494];
    assign line_data_495 = line_data[495];
    assign line_data_496 = line_data[496];
    assign line_data_497 = line_data[497];
    assign line_data_498 = line_data[498];
    assign line_data_499 = line_data[499];
    assign line_data_500 = line_data[500];
    assign line_data_501 = line_data[501];
    assign line_data_502 = line_data[502];
    assign line_data_503 = line_data[503];
    assign line_data_504 = line_data[504];
    assign line_data_505 = line_data[505];
    assign line_data_506 = line_data[506];
    assign line_data_507 = line_data[507];
    assign line_data_508 = line_data[508];
    assign line_data_509 = line_data[509];
    assign line_data_510 = line_data[510];
    assign line_data_511 = line_data[511];
    assign line_data_512 = line_data[512];
    assign line_data_513 = line_data[513];
    assign line_data_514 = line_data[514];
    assign line_data_515 = line_data[515];
    assign line_data_516 = line_data[516];
    assign line_data_517 = line_data[517];
    assign line_data_518 = line_data[518];
    assign line_data_519 = line_data[519];
    assign line_data_520 = line_data[520];
    assign line_data_521 = line_data[521];
    assign line_data_522 = line_data[522];
    assign line_data_523 = line_data[523];
    assign line_data_524 = line_data[524];
    assign line_data_525 = line_data[525];
    assign line_data_526 = line_data[526];
    assign line_data_527 = line_data[527];
    assign line_data_528 = line_data[528];
    assign line_data_529 = line_data[529];
    assign line_data_530 = line_data[530];
    assign line_data_531 = line_data[531];
    assign line_data_532 = line_data[532];
    assign line_data_533 = line_data[533];
    assign line_data_534 = line_data[534];
    assign line_data_535 = line_data[535];
    assign line_data_536 = line_data[536];
    assign line_data_537 = line_data[537];
    assign line_data_538 = line_data[538];
    assign line_data_539 = line_data[539];
    assign line_data_540 = line_data[540];
    assign line_data_541 = line_data[541];
    assign line_data_542 = line_data[542];
    assign line_data_543 = line_data[543];
    assign line_data_544 = line_data[544];
    assign line_data_545 = line_data[545];
    assign line_data_546 = line_data[546];
    assign line_data_547 = line_data[547];
    assign line_data_548 = line_data[548];
    assign line_data_549 = line_data[549];
    assign line_data_550 = line_data[550];
    assign line_data_551 = line_data[551];
    assign line_data_552 = line_data[552];
    assign line_data_553 = line_data[553];
    assign line_data_554 = line_data[554];
    assign line_data_555 = line_data[555];
    assign line_data_556 = line_data[556];
    assign line_data_557 = line_data[557];
    assign line_data_558 = line_data[558];
    assign line_data_559 = line_data[559];
    assign line_data_560 = line_data[560];
    assign line_data_561 = line_data[561];
    assign line_data_562 = line_data[562];
    assign line_data_563 = line_data[563];
    assign line_data_564 = line_data[564];
    assign line_data_565 = line_data[565];
    assign line_data_566 = line_data[566];
    assign line_data_567 = line_data[567];
    assign line_data_568 = line_data[568];
    assign line_data_569 = line_data[569];
    assign line_data_570 = line_data[570];
    assign line_data_571 = line_data[571];
    assign line_data_572 = line_data[572];
    assign line_data_573 = line_data[573];
    assign line_data_574 = line_data[574];
    assign line_data_575 = line_data[575];
    assign line_data_576 = line_data[576];
    assign line_data_577 = line_data[577];
    assign line_data_578 = line_data[578];
    assign line_data_579 = line_data[579];
    assign line_data_580 = line_data[580];
    assign line_data_581 = line_data[581];
    assign line_data_582 = line_data[582];
    assign line_data_583 = line_data[583];
    assign line_data_584 = line_data[584];
    assign line_data_585 = line_data[585];
    assign line_data_586 = line_data[586];
    assign line_data_587 = line_data[587];
    assign line_data_588 = line_data[588];
    assign line_data_589 = line_data[589];
    assign line_data_590 = line_data[590];
    assign line_data_591 = line_data[591];
    assign line_data_592 = line_data[592];
    assign line_data_593 = line_data[593];
    assign line_data_594 = line_data[594];
    assign line_data_595 = line_data[595];
    assign line_data_596 = line_data[596];
    assign line_data_597 = line_data[597];
    assign line_data_598 = line_data[598];
    assign line_data_599 = line_data[599];
    assign line_data_600 = line_data[600];
    assign line_data_601 = line_data[601];
    assign line_data_602 = line_data[602];
    assign line_data_603 = line_data[603];
    assign line_data_604 = line_data[604];
    assign line_data_605 = line_data[605];
    assign line_data_606 = line_data[606];
    assign line_data_607 = line_data[607];
    assign line_data_608 = line_data[608];
    assign line_data_609 = line_data[609];
    assign line_data_610 = line_data[610];
    assign line_data_611 = line_data[611];
    assign line_data_612 = line_data[612];
    assign line_data_613 = line_data[613];
    assign line_data_614 = line_data[614];
    assign line_data_615 = line_data[615];
    assign line_data_616 = line_data[616];
    assign line_data_617 = line_data[617];
    assign line_data_618 = line_data[618];
    assign line_data_619 = line_data[619];
    assign line_data_620 = line_data[620];
    assign line_data_621 = line_data[621];
    assign line_data_622 = line_data[622];
    assign line_data_623 = line_data[623];
    assign line_data_624 = line_data[624];
    assign line_data_625 = line_data[625];
    assign line_data_626 = line_data[626];
    assign line_data_627 = line_data[627];
    assign line_data_628 = line_data[628];
    assign line_data_629 = line_data[629];
    assign line_data_630 = line_data[630];
    assign line_data_631 = line_data[631];
    assign line_data_632 = line_data[632];
    assign line_data_633 = line_data[633];
    assign line_data_634 = line_data[634];
    assign line_data_635 = line_data[635];
    assign line_data_636 = line_data[636];
    assign line_data_637 = line_data[637];
    assign line_data_638 = line_data[638];
    assign line_data_639 = line_data[639];
    assign line_data_640 = line_data[640];
    assign line_data_641 = line_data[641];
    assign line_data_642 = line_data[642];
    assign line_data_643 = line_data[643];
    assign line_data_644 = line_data[644];
    assign line_data_645 = line_data[645];
    assign line_data_646 = line_data[646];
    assign line_data_647 = line_data[647];
    assign line_data_648 = line_data[648];
    assign line_data_649 = line_data[649];
    assign line_data_650 = line_data[650];
    assign line_data_651 = line_data[651];
    assign line_data_652 = line_data[652];
    assign line_data_653 = line_data[653];
    assign line_data_654 = line_data[654];
    assign line_data_655 = line_data[655];
    assign line_data_656 = line_data[656];
    assign line_data_657 = line_data[657];
    assign line_data_658 = line_data[658];
    assign line_data_659 = line_data[659];
    assign line_data_660 = line_data[660];
    assign line_data_661 = line_data[661];
    assign line_data_662 = line_data[662];
    assign line_data_663 = line_data[663];
    assign line_data_664 = line_data[664];
    assign line_data_665 = line_data[665];
    assign line_data_666 = line_data[666];
    assign line_data_667 = line_data[667];
    assign line_data_668 = line_data[668];
    assign line_data_669 = line_data[669];
    assign line_data_670 = line_data[670];
    assign line_data_671 = line_data[671];
    assign line_data_672 = line_data[672];
    assign line_data_673 = line_data[673];
    assign line_data_674 = line_data[674];
    assign line_data_675 = line_data[675];
    assign line_data_676 = line_data[676];
    assign line_data_677 = line_data[677];
    assign line_data_678 = line_data[678];
    assign line_data_679 = line_data[679];
    assign line_data_680 = line_data[680];
    assign line_data_681 = line_data[681];
    assign line_data_682 = line_data[682];
    assign line_data_683 = line_data[683];
    assign line_data_684 = line_data[684];
    assign line_data_685 = line_data[685];
    assign line_data_686 = line_data[686];
    assign line_data_687 = line_data[687];
    assign line_data_688 = line_data[688];
    assign line_data_689 = line_data[689];
    assign line_data_690 = line_data[690];
    assign line_data_691 = line_data[691];
    assign line_data_692 = line_data[692];
    assign line_data_693 = line_data[693];
    assign line_data_694 = line_data[694];
    assign line_data_695 = line_data[695];
    assign line_data_696 = line_data[696];
    assign line_data_697 = line_data[697];
    assign line_data_698 = line_data[698];
    assign line_data_699 = line_data[699];
    assign line_data_700 = line_data[700];
    assign line_data_701 = line_data[701];
    assign line_data_702 = line_data[702];
    assign line_data_703 = line_data[703];
    assign line_data_704 = line_data[704];
    assign line_data_705 = line_data[705];
    assign line_data_706 = line_data[706];
    assign line_data_707 = line_data[707];
    assign line_data_708 = line_data[708];
    assign line_data_709 = line_data[709];
    assign line_data_710 = line_data[710];
    assign line_data_711 = line_data[711];
    assign line_data_712 = line_data[712];
    assign line_data_713 = line_data[713];
    assign line_data_714 = line_data[714];
    assign line_data_715 = line_data[715];
    assign line_data_716 = line_data[716];
    assign line_data_717 = line_data[717];
    assign line_data_718 = line_data[718];
    assign line_data_719 = line_data[719];
    assign line_data_720 = line_data[720];
    assign line_data_721 = line_data[721];
    assign line_data_722 = line_data[722];
    assign line_data_723 = line_data[723];
    assign line_data_724 = line_data[724];
    assign line_data_725 = line_data[725];
    assign line_data_726 = line_data[726];
    assign line_data_727 = line_data[727];
    assign line_data_728 = line_data[728];
    assign line_data_729 = line_data[729];
    assign line_data_730 = line_data[730];
    assign line_data_731 = line_data[731];
    assign line_data_732 = line_data[732];
    assign line_data_733 = line_data[733];
    assign line_data_734 = line_data[734];
    assign line_data_735 = line_data[735];
    assign line_data_736 = line_data[736];
    assign line_data_737 = line_data[737];
    assign line_data_738 = line_data[738];
    assign line_data_739 = line_data[739];
    assign line_data_740 = line_data[740];
    assign line_data_741 = line_data[741];
    assign line_data_742 = line_data[742];
    assign line_data_743 = line_data[743];
    assign line_data_744 = line_data[744];
    assign line_data_745 = line_data[745];
    assign line_data_746 = line_data[746];
    assign line_data_747 = line_data[747];
    assign line_data_748 = line_data[748];
    assign line_data_749 = line_data[749];
    assign line_data_750 = line_data[750];
    assign line_data_751 = line_data[751];
    assign line_data_752 = line_data[752];
    assign line_data_753 = line_data[753];
    assign line_data_754 = line_data[754];
    assign line_data_755 = line_data[755];
    assign line_data_756 = line_data[756];
    assign line_data_757 = line_data[757];
    assign line_data_758 = line_data[758];
    assign line_data_759 = line_data[759];
    assign line_data_760 = line_data[760];
    assign line_data_761 = line_data[761];
    assign line_data_762 = line_data[762];
    assign line_data_763 = line_data[763];
    assign line_data_764 = line_data[764];
    assign line_data_765 = line_data[765];
    assign line_data_766 = line_data[766];
    assign line_data_767 = line_data[767];
    assign line_data_768 = line_data[768];
    assign line_data_769 = line_data[769];
    assign line_data_770 = line_data[770];
    assign line_data_771 = line_data[771];
    assign line_data_772 = line_data[772];
    assign line_data_773 = line_data[773];
    assign line_data_774 = line_data[774];
    assign line_data_775 = line_data[775];
    assign line_data_776 = line_data[776];
    assign line_data_777 = line_data[777];
    assign line_data_778 = line_data[778];
    assign line_data_779 = line_data[779];
    assign line_data_780 = line_data[780];
    assign line_data_781 = line_data[781];
    assign line_data_782 = line_data[782];
    assign line_data_783 = line_data[783];
    assign line_data_784 = line_data[784];
    assign line_data_785 = line_data[785];
    assign line_data_786 = line_data[786];
    assign line_data_787 = line_data[787];
    assign line_data_788 = line_data[788];
    assign line_data_789 = line_data[789];
    assign line_data_790 = line_data[790];
    assign line_data_791 = line_data[791];
    assign line_data_792 = line_data[792];
    assign line_data_793 = line_data[793];
    assign line_data_794 = line_data[794];
    assign line_data_795 = line_data[795];
    assign line_data_796 = line_data[796];
    assign line_data_797 = line_data[797];
    assign line_data_798 = line_data[798];
    assign line_data_799 = line_data[799];
    assign line_data_800 = line_data[800];
    assign line_data_801 = line_data[801];
    assign line_data_802 = line_data[802];
    assign line_data_803 = line_data[803];
    assign line_data_804 = line_data[804];
    assign line_data_805 = line_data[805];
    assign line_data_806 = line_data[806];
    assign line_data_807 = line_data[807];
    assign line_data_808 = line_data[808];
    assign line_data_809 = line_data[809];
    assign line_data_810 = line_data[810];
    assign line_data_811 = line_data[811];
    assign line_data_812 = line_data[812];
    assign line_data_813 = line_data[813];
    assign line_data_814 = line_data[814];
    assign line_data_815 = line_data[815];
    assign line_data_816 = line_data[816];
    assign line_data_817 = line_data[817];
    assign line_data_818 = line_data[818];
    assign line_data_819 = line_data[819];
    assign line_data_820 = line_data[820];
    assign line_data_821 = line_data[821];
    assign line_data_822 = line_data[822];
    assign line_data_823 = line_data[823];
    assign line_data_824 = line_data[824];
    assign line_data_825 = line_data[825];
    assign line_data_826 = line_data[826];
    assign line_data_827 = line_data[827];
    assign line_data_828 = line_data[828];
    assign line_data_829 = line_data[829];
    assign line_data_830 = line_data[830];
    assign line_data_831 = line_data[831];
    assign line_data_832 = line_data[832];
    assign line_data_833 = line_data[833];
    assign line_data_834 = line_data[834];
    assign line_data_835 = line_data[835];
    assign line_data_836 = line_data[836];
    assign line_data_837 = line_data[837];
    assign line_data_838 = line_data[838];
    assign line_data_839 = line_data[839];
    assign line_data_840 = line_data[840];
    assign line_data_841 = line_data[841];
    assign line_data_842 = line_data[842];
    assign line_data_843 = line_data[843];
    assign line_data_844 = line_data[844];
    assign line_data_845 = line_data[845];
    assign line_data_846 = line_data[846];
    assign line_data_847 = line_data[847];
    assign line_data_848 = line_data[848];
    assign line_data_849 = line_data[849];
    assign line_data_850 = line_data[850];
    assign line_data_851 = line_data[851];
    assign line_data_852 = line_data[852];
    assign line_data_853 = line_data[853];
    assign line_data_854 = line_data[854];
    assign line_data_855 = line_data[855];
    assign line_data_856 = line_data[856];
    assign line_data_857 = line_data[857];
    assign line_data_858 = line_data[858];
    assign line_data_859 = line_data[859];
    assign line_data_860 = line_data[860];
    assign line_data_861 = line_data[861];
    assign line_data_862 = line_data[862];
    assign line_data_863 = line_data[863];
    assign line_data_864 = line_data[864];
    assign line_data_865 = line_data[865];
    assign line_data_866 = line_data[866];
    assign line_data_867 = line_data[867];
    assign line_data_868 = line_data[868];
    assign line_data_869 = line_data[869];
    assign line_data_870 = line_data[870];
    assign line_data_871 = line_data[871];
    assign line_data_872 = line_data[872];
    assign line_data_873 = line_data[873];
    assign line_data_874 = line_data[874];
    assign line_data_875 = line_data[875];
    assign line_data_876 = line_data[876];
    assign line_data_877 = line_data[877];
    assign line_data_878 = line_data[878];
    assign line_data_879 = line_data[879];
    assign line_data_880 = line_data[880];
    assign line_data_881 = line_data[881];
    assign line_data_882 = line_data[882];
    assign line_data_883 = line_data[883];
    assign line_data_884 = line_data[884];
    assign line_data_885 = line_data[885];
    assign line_data_886 = line_data[886];
    assign line_data_887 = line_data[887];
    assign line_data_888 = line_data[888];
    assign line_data_889 = line_data[889];
    assign line_data_890 = line_data[890];
    assign line_data_891 = line_data[891];
    assign line_data_892 = line_data[892];
    assign line_data_893 = line_data[893];
    assign line_data_894 = line_data[894];
    assign line_data_895 = line_data[895];
    assign line_data_896 = line_data[896];
    assign line_data_897 = line_data[897];
    assign line_data_898 = line_data[898];
    assign line_data_899 = line_data[899];
    assign line_data_900 = line_data[900];
    assign line_data_901 = line_data[901];
    assign line_data_902 = line_data[902];
    assign line_data_903 = line_data[903];
    assign line_data_904 = line_data[904];
    assign line_data_905 = line_data[905];
    assign line_data_906 = line_data[906];
    assign line_data_907 = line_data[907];
    assign line_data_908 = line_data[908];
    assign line_data_909 = line_data[909];
    assign line_data_910 = line_data[910];
    assign line_data_911 = line_data[911];
    assign line_data_912 = line_data[912];
    assign line_data_913 = line_data[913];
    assign line_data_914 = line_data[914];
    assign line_data_915 = line_data[915];
    assign line_data_916 = line_data[916];
    assign line_data_917 = line_data[917];
    assign line_data_918 = line_data[918];
    assign line_data_919 = line_data[919];
    assign line_data_920 = line_data[920];
    assign line_data_921 = line_data[921];
    assign line_data_922 = line_data[922];
    assign line_data_923 = line_data[923];
    assign line_data_924 = line_data[924];
    assign line_data_925 = line_data[925];
    assign line_data_926 = line_data[926];
    assign line_data_927 = line_data[927];
    assign line_data_928 = line_data[928];
    assign line_data_929 = line_data[929];
    assign line_data_930 = line_data[930];
    assign line_data_931 = line_data[931];
    assign line_data_932 = line_data[932];
    assign line_data_933 = line_data[933];
    assign line_data_934 = line_data[934];
    assign line_data_935 = line_data[935];
    assign line_data_936 = line_data[936];
    assign line_data_937 = line_data[937];
    assign line_data_938 = line_data[938];
    assign line_data_939 = line_data[939];
    assign line_data_940 = line_data[940];
    assign line_data_941 = line_data[941];
    assign line_data_942 = line_data[942];
    assign line_data_943 = line_data[943];
    assign line_data_944 = line_data[944];
    assign line_data_945 = line_data[945];
    assign line_data_946 = line_data[946];
    assign line_data_947 = line_data[947];
    assign line_data_948 = line_data[948];
    assign line_data_949 = line_data[949];
    assign line_data_950 = line_data[950];
    assign line_data_951 = line_data[951];
    assign line_data_952 = line_data[952];
    assign line_data_953 = line_data[953];
    assign line_data_954 = line_data[954];
    assign line_data_955 = line_data[955];
    assign line_data_956 = line_data[956];
    assign line_data_957 = line_data[957];
    assign line_data_958 = line_data[958];
    assign line_data_959 = line_data[959];
    assign line_data_960 = line_data[960];
    assign line_data_961 = line_data[961];
    assign line_data_962 = line_data[962];
    assign line_data_963 = line_data[963];
    assign line_data_964 = line_data[964];
    assign line_data_965 = line_data[965];
    assign line_data_966 = line_data[966];
    assign line_data_967 = line_data[967];
    assign line_data_968 = line_data[968];
    assign line_data_969 = line_data[969];
    assign line_data_970 = line_data[970];
    assign line_data_971 = line_data[971];
    assign line_data_972 = line_data[972];
    assign line_data_973 = line_data[973];
    assign line_data_974 = line_data[974];
    assign line_data_975 = line_data[975];
    assign line_data_976 = line_data[976];
    assign line_data_977 = line_data[977];
    assign line_data_978 = line_data[978];
    assign line_data_979 = line_data[979];
    assign line_data_980 = line_data[980];
    assign line_data_981 = line_data[981];
    assign line_data_982 = line_data[982];
    assign line_data_983 = line_data[983];
    assign line_data_984 = line_data[984];
    assign line_data_985 = line_data[985];
    assign line_data_986 = line_data[986];
    assign line_data_987 = line_data[987];
    assign line_data_988 = line_data[988];
    assign line_data_989 = line_data[989];
    assign line_data_990 = line_data[990];
    assign line_data_991 = line_data[991];
    assign line_data_992 = line_data[992];
    assign line_data_993 = line_data[993];
    assign line_data_994 = line_data[994];
    assign line_data_995 = line_data[995];
    assign line_data_996 = line_data[996];
    assign line_data_997 = line_data[997];
    assign line_data_998 = line_data[998];
    assign line_data_999 = line_data[999];
    assign line_data_1000 = line_data[1000];
    assign line_data_1001 = line_data[1001];
    assign line_data_1002 = line_data[1002];
    assign line_data_1003 = line_data[1003];
    assign line_data_1004 = line_data[1004];
    assign line_data_1005 = line_data[1005];
    assign line_data_1006 = line_data[1006];
    assign line_data_1007 = line_data[1007];
    assign line_data_1008 = line_data[1008];
    assign line_data_1009 = line_data[1009];
    assign line_data_1010 = line_data[1010];
    assign line_data_1011 = line_data[1011];
    assign line_data_1012 = line_data[1012];
    assign line_data_1013 = line_data[1013];
    assign line_data_1014 = line_data[1014];
    assign line_data_1015 = line_data[1015];
    assign line_data_1016 = line_data[1016];
    assign line_data_1017 = line_data[1017];
    assign line_data_1018 = line_data[1018];
    assign line_data_1019 = line_data[1019];
    assign line_data_1020 = line_data[1020];
    assign line_data_1021 = line_data[1021];
    assign line_data_1022 = line_data[1022];
    assign line_data_1023 = line_data[1023];
    
       
    
       always @(*) begin
           softmax_read_FP16_matrix(en, line_num, line_data); 
       end
    
endmodule

