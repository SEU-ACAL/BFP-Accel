module tb(
  input   clock,
  input   reset
);
endmodule
